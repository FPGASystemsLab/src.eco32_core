//==============================================================================================
//    Main contributors
//      - Adam Luczak         <mailto:adam.luczak@outlook.com>
//==============================================================================================
`default_nettype none
//----------------------------------------------------------------------------------------------
`timescale 1ns / 1ns                            
//==============================================================================================
module eco32_core_mpu_erx 
(
 input  wire         clk,
 input  wire         rst,

 input  wire   [8:0] wr_bus,

 input  wire         rd_tid,
 input  wire   [3:0] rd_addr,
 output wire  [63:0] rd_data
);
//==============================================================================================
//  params
//==============================================================================================
parameter               FORCE_RST   =     0;
//==============================================================================================
// variables
//==============================================================================================
reg     [63:0]  erx [31:0]; 
reg     [71:0]  wr_buff; // 64 + {1(tid),4(addr)}
reg             wr_tag; 
//==============================================================================================
// deserialiser
//==============================================================================================
always@(posedge clk or posedge rst)
 if(rst)    wr_buff                 <=                                                      'd0;        
 else       wr_buff                 <=                              {wr_bus[7:0],wr_buff[71:8]};        
//----------------------------------------------------------------------------------------------         
always@(posedge clk or posedge rst)                                                                          
 if(rst)    wr_tag                  <=                                                      'd0;        
 else       wr_tag                  <=                                                wr_bus[8];        
//==============================================================================================
wire        wr_ena                   =                                                   wr_tag;
wire        wr_tid                   =                                           wr_buff[   68];
wire  [3:0] wr_addr                  =                                           wr_buff[67:64];
wire [63:0] wr_data                  =                                           wr_buff[63: 0];
//----------------------------------------------------------------------------------------------
always@(posedge clk)
 if(wr_ena) erx[{wr_tid,wr_addr}]  <=                                                   wr_data;
//----------------------------------------------------------------------------------------------
assign      rd_data                 =                                     erx[{rd_tid,rd_addr}];
//==============================================================================================
endmodule                                                                                   
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            