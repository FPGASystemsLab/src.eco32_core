//=============================================================================
//    Main contributors
//      - Adam Luczak         <mailto:adam.luczak@outlook.com>
//=============================================================================
`default_nettype none
//-----------------------------------------------------------------------------
`timescale 1ns / 1ns                            
//=============================================================================
module eco32_core_idu_rfu_reg 
(                        
 input  wire            clk,

 input  wire     [4:0]  i_addr,

 input  wire            w_ena,     
 input  wire     [3:0]  w_ben,
 input  wire     [4:0]  w_addr,
 input  wire    [31:0]  w_data,
 
 output wire    [31:0]  o_data
);                             
//=============================================================================
// variable
//=============================================================================
reg     [7:0]   mem_b0  [0:31]; /* synthesis ramstyle = "distributed" */
reg     [7:0]   mem_b1  [0:31]; /* synthesis ramstyle = "distributed" */ 
reg     [7:0]   mem_b2  [0:31]; /* synthesis ramstyle = "distributed" */
reg     [7:0]   mem_b3  [0:31]; /* synthesis ramstyle = "distributed" */
//-----------------------------------------------------------------------------
wire            wen0    =   w_ena & w_ben[0];
wire            wen1    =   w_ena & w_ben[1];
wire            wen2    =   w_ena & w_ben[2];
wire            wen3    =   w_ena & w_ben[3];
//=============================================================================
// memory
//=============================================================================
always@(posedge clk) if(wen0) mem_b0[w_addr] <= w_data[7:0];
//-----------------------------------------------------------------------------
assign  o_data[7:0] = mem_b0[i_addr];
//=============================================================================
always@(posedge clk) if(wen1) mem_b1[w_addr] <= w_data[15:8];
//-----------------------------------------------------------------------------
assign  o_data[15:8] = mem_b1[i_addr];
//=============================================================================
always@(posedge clk) if(wen2) mem_b2[w_addr] <= w_data[23:16];
//-----------------------------------------------------------------------------
assign  o_data[23:16] = mem_b2[i_addr];
//=============================================================================
always@(posedge clk) if(wen3) mem_b3[w_addr] <= w_data[31:24];
//-----------------------------------------------------------------------------
assign  o_data[31:24] = mem_b3[i_addr];
//=============================================================================
endmodule