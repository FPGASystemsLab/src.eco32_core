//==============================================================================================
//    Main contributors
//      - Adam Luczak         <mailto:adam.luczak@outlook.com>
//==============================================================================================
`default_nettype none
//----------------------------------------------------------------------------------------------
`timescale 1ns / 1ns                            
//==============================================================================================
module eco32_core_mpu_crx 
(
 input  wire         clk,
 input  wire         rst,

 input  wire         i_tid,
 input  wire   [4:0] i_addr,
 input  wire         i_wra,     
 input  wire  [31:0] i_cra,
 input  wire         i_wrb,     
 input  wire         i_wri,     
 input  wire  [31:0] i_crb,     

 output wire  [31:0] o_cra,
 output wire  [31:0] o_crb,       
 
 output wire   [5:0] sys_asid,     
 output wire   [1:0] sys_trace_ena,
 output wire   [1:0] sys_event_ena
);
//==============================================================================================
// variables
//==============================================================================================
reg     [31:0]  cra [63:0]; 
reg     [30:0]  crx [63:0];
reg             cri [63:0];
//----------------------------------------------------------------------------------------------
reg     [5:0]   scf_asid_a;
reg     [5:0]   scf_asid_b;
//----------------------------------------------------------------------------------------------
reg             scf_tid;
//----------------------------------------------------------------------------------------------
reg             scf_event_enable_th0;
reg             scf_event_enable_th1;
//----------------------------------------------------------------------------------------------
reg             scf_trace_enable_th0;
reg             scf_trace_enable_th1;
//============================================================================================== 
// cra regs
//============================================================================================== 
always@(posedge clk)
 if(i_wra)          cra [{i_tid,i_addr}] <=                                                i_cra;
//----------------------------------------------------------------------------------------------
wire    [31:0]      cra_out      =                                         cra [{i_tid,i_addr}];
//============================================================================================== 
// crb regs
//============================================================================================== 
always@(posedge clk)
 if(i_wrb)          crx [{i_tid,i_addr}] <=                                         i_crb[31:1];
//----------------------------------------------------------------------------------------------
always@(posedge clk)
 if(i_wri)          cri [{i_tid,i_addr}] <=                                            i_crb[0];
//----------------------------------------------------------------------------------------------
wire    [31:0]      crb_out          =              {crx [{i_tid,i_addr}],cri [{i_tid,i_addr}]};                                     
//============================================================================================== 
// output 
//============================================================================================== 
assign              o_cra            =                                                  cra_out;
assign              o_crb            =                                                  crb_out;
//==============================================================================================
// system control flags
//==============================================================================================
// address space [5:0]
//----------------------------------------------------------------------------------------------
wire            f_asid           =                                                i_addr==5'd08;
wire            f_trace_enable0  =                                 i_tid==1'b0 && i_addr==5'd10;
wire            f_trace_enable1  =                                 i_tid==1'b1 && i_addr==5'd10;
wire            f_event_enable0  =                                 i_tid==1'b0 && i_addr==5'd14;
wire            f_event_enable1  =                                 i_tid==1'b1 && i_addr==5'd14;
//==============================================================================================
// tid buffer
//==============================================================================================
always@(posedge clk or posedge rst)
 if(rst)                                scf_tid             <=                              'd0;    
 else                                   scf_tid             <=                            i_tid;    
//==============================================================================================
// assid 
//==============================================================================================
always@(posedge clk or posedge rst)
 if(rst)                                scf_asid_a          <=                              'd0;
 else if(i_wra && f_asid)               scf_asid_a          <=                       i_crb[5:0];
 else                                   scf_asid_a          <=                       scf_asid_b;
//---------------------------------------------------------------------------------------------
always@(posedge clk or posedge rst)
 if(rst)                                scf_asid_b          <=                              'd0;    
 else                                   scf_asid_b          <=                       scf_asid_a;    
//---------------------------------------------------------------------------------------------
assign                                  sys_asid             =                       scf_asid_a;
//==============================================================================================
// event enable
//==============================================================================================
always@(posedge clk or posedge rst)
 if(rst)                                scf_event_enable_th0<=                              'd0;  
 else if(i_wri && f_event_enable0)      scf_event_enable_th0<=                         i_crb[0];
//----------------------------------------------------------------------------------------------
assign                                  sys_event_ena[0]     =             scf_event_enable_th0;
//----------------------------------------------------------------------------------------------
always@(posedge clk or posedge rst)
 if(rst)                                scf_event_enable_th1<=                              'd0;  
 else if(i_wri && f_event_enable1)      scf_event_enable_th1<=                         i_crb[0];                         
//----------------------------------------------------------------------------------------------
assign                                  sys_event_ena[1]     =             scf_event_enable_th1;
//==============================================================================================
always@(posedge clk or posedge rst)
 if(rst)                                scf_trace_enable_th0<=                              'd0;    
 else if(i_wrb && f_trace_enable0)      scf_trace_enable_th0<=                         i_crb[0];
//----------------------------------------------------------------------------------------------
assign                                  sys_trace_ena[0]     =             scf_trace_enable_th0;
//----------------------------------------------------------------------------------------------
always@(posedge clk or posedge rst)
 if(rst)                                scf_trace_enable_th1<=                              'd0;
 else if(i_wrb && f_trace_enable1)      scf_trace_enable_th1<=                         i_crb[0];
//----------------------------------------------------------------------------------------------
assign                                  sys_trace_ena[1]     =             scf_trace_enable_th1;
//==============================================================================================
endmodule                                                                                   
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            