//==============================================================================================
//    Main contributors
//      - Adam Luczak         <mailto:adam.luczak@outlook.com>
//==============================================================================================
`default_nettype none
//----------------------------------------------------------------------------------------------
`timescale 1ns / 1ns                            
//==============================================================================================
module eco32_core_mpu_cfr 
(
 input  wire         clk,
 input  wire         rst,

 input  wire         ia_wen,     
 input  wire  [15:0] ia_flags,     
 
 input  wire         ib_wen,     
 input  wire  [15:0] ib_flags,     

 output wire  [15:0] o_flags,
 
 output wire         dbg_stb,
 output wire   [6:0] dbg_flags
);
//==============================================================================================
// variables
//==============================================================================================
reg        b1_flags_change; 
reg [15:0] b1_flags; 
reg [15:0] a2_flags; 
//==============================================================================================
// flags for th 0
//==============================================================================================
always@(posedge clk or posedge rst)
 if(rst)            b1_flags        <=                                                    16'd0;
 else if(ia_wen)    b1_flags        <=                                                 ia_flags;
 else if(ib_wen)    b1_flags        <=                                                 ib_flags;
 else               b1_flags        <=                                                 a2_flags;
//----------------------------------------------------------------------------------------------
always@(posedge clk or posedge rst)
 if(rst)            b1_flags_change <=                                                     1'd0;
 else if(ia_wen)    b1_flags_change <=                                                     1'd1;
 else if(ib_wen)    b1_flags_change <=                                                     1'd1;
 else               b1_flags_change <=                                                     1'd0;
//==============================================================================================
// b3
//==============================================================================================
always@(posedge clk or posedge rst)
 if(rst)            a2_flags        <=                                                    12'd0;
 else               a2_flags        <=                                                 b1_flags;
//==============================================================================================
assign              o_flags          =                                                 b1_flags;
//==============================================================================================    
// debug
//==============================================================================================    
assign              dbg_stb          =                                          b1_flags_change;
assign              dbg_flags        =                            {b1_flags[9:7],b1_flags[3:0]};
//==============================================================================================    
endmodule                                                                                   
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            
                                                                                            