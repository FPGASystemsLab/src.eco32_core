//=============================================================================
//    Main contributors
//      - Adam Luczak         <mailto:adam.luczak@outlook.com>
//=============================================================================
`default_nettype none
//-----------------------------------------------------------------------------
`timescale 1ns / 1ns                            
//=============================================================================
module eco32_core_idu_rfu_tag 
(                        
 input  wire            clk,

 input  wire     [4:0]  i_addr,

 input  wire            w_ena,     
 input  wire     [4:0]  w_addr,     
 input  wire            w_tag,    
 
 output wire            o_tag
);                             
//=============================================================================
// variable
//=============================================================================
reg     [31:0]  mem; /* synthesis ramstyle = "distributed" */
//=============================================================================
// memory
//=============================================================================
always@(posedge clk) if(w_ena) mem[w_addr] <= w_tag;
//-----------------------------------------------------------------------------          
assign  o_tag = mem[i_addr];                                                          
//=============================================================================
endmodule