//==============================================================================================
//    Main contributors
//      - Adam Luczak         <mailto:adam.luczak@outlook.com>
//==============================================================================================
`default_nettype none
//----------------------------------------------------------------------------------------------
`timescale 1ns / 1ns                            
//==============================================================================================
// hierarchy:
// processor core (TOP)
// + instruction fetch 
//   + instruction cache way 
//     + instruction cache memory
//==============================================================================================
module eco32_core_ifu_icu_way_mem 
# // parameters
(
parameter [5:0]  PAGE_ADDR_WIDTH  =  6'h5
)
// ports
(
input  wire                             clk,

input  wire                             i_tid,
input  wire  [PAGE_ADDR_WIDTH-1:0]  i_page,
input  wire                    [2:0]    i_offset,     

input  wire                             wr_ena,
input  wire                             wr_tid,
input  wire  [PAGE_ADDR_WIDTH-1:0]  wr_page,
input  wire                    [2:0]    wr_offset,
input  wire                   [71:0]    wr_data,
 
output wire                   [71:0]    o_data
);                             
//==============================================================================================
// parameters
//==============================================================================================
localparam          _A                  =                             (PAGE_ADDR_WIDTH + 1 + 3);
localparam          _P                  =                             (PAGE_ADDR_WIDTH        );
localparam          _T                  =                          1<<(PAGE_ADDR_WIDTH + 1 + 3);       
//==============================================================================================
// variables
//==============================================================================================
(*ramstyle="no_rw_check"*) reg     [  71:0] mem [_T-1:0];
                           reg     [_A-1:0] mem_ptr;    
                           wire    [_A-1:0] wr_addr;
                           wire    [_A-1:0] rd_addr;
                           wire    [  71:0] rd_data;    
//==============================================================================================
// memory
//==============================================================================================
assign  wr_addr     =                                                {wr_page,wr_tid,wr_offset};
assign  rd_addr     =                                                {  i_page,i_tid, i_offset};
//----------------------------------------------------------------------------------------------
always@(posedge clk)
    begin
        if(wr_ena)  mem[wr_addr]    <= wr_data;
        mem_ptr                     <= rd_addr;
    end
//----------------------------------------------------------------------------------------------
assign  rd_data     =                                                              mem[mem_ptr];
//==============================================================================================
assign  o_data      =                                                                   rd_data;
//==============================================================================================
endmodule